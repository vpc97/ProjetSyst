`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    08:52:25 05/17/2018 
// Design Name: 
// Module Name:    bancregistres 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module bancregistres(
    input @A,
    input @B,
    input RST,
    input CLK,
    output QA,
    output QB,
    input @W,
    input W,
    input DATA
    );


endmodule
